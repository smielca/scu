module main

import scu

pub struct Button {
	scu.Node
pub mut:
    button_text string
}
